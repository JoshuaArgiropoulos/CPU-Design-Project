module RAM_Reg(input Data_Signal[31:0], input Read, input Write, input Address_Signal[31:0], output BusMuxIn)
  
