`timescale 1ns/10ps
module DP_Branch_TB;

reg [31:0] enable, busSelect, inPort, MDataIn;
reg clk, clr, MD_Read, Gra, Grb, Grc, Rin, Rout, BAout, WriteRAM, ReadRAM;//, IncPC;
reg [4:0] Control_Signals;
wire [31:0] busMuxOut, r1, r2, r3, mdr, zhi, zlo, pc, ir;//, hi, lo, temp;
//wire [63:0] temp;

parameter Default = 4'b0000, Reg_load1a = 4'b0001, Reg_load1b = 4'b0010, Reg_load2a = 4'b0011, 
			 Reg_load2b = 4'b0100, Reg_load3a = 4'b0101, Reg_load3b = 4'b0110, T0 = 4'b0111, 
			 T1 = 4'b1000, T2 = 4'b1001, T3 = 4'b1010, T4 = 4'b1011, T5 = 4'b1100, T6 = 4'b1101, T7 = 4'b1110;
reg [3:0] Present_state = Default;

	 

datapath DUT(enable, busSelect, inPort, /*MDataIn,*/ clk, clr, MD_Read, Gra, Grb, Grc, Rin, Rout, BAout, WriteRAM, ReadRAM, Control_Signals, busMuxOut, r1, r2, r3, mdr, zhi, zlo, pc, ir);//, hi, lo, temp); 



initial begin

clk = 0;
forever #10 clk = ~clk;

end

always @(posedge clk) begin
	case(Present_state)
		Default : Present_state = Reg_load1a;
		Reg_load1a :#40 Present_state = Reg_load1b;
		Reg_load1b :#40 Present_state = Reg_load2a;
		Reg_load2a :#40 Present_state = Reg_load2b;
		Reg_load2b :#40 Present_state = Reg_load3a;
		Reg_load3a :#40 Present_state = Reg_load3b;
		Reg_load3b :#40 Present_state = T0;
		T0 :#40 Present_state = T1;
		T1 :#40 Present_state = T2;
		T2 :#40 Present_state = T3;
		T3 :#40 Present_state = T4;
		T4 :#40 Present_state = T5;
		T5 :#40 Present_state = T6;
		T6 :#40 Present_state = T7;
	endcase
end

always @(Present_state) begin

	case(Present_state)
	
	
		Default: begin
								busSelect <= 32'b0;
								enable <= 32'b0;
								MD_Read <= 0;
								Control_Signals <= 4'b0;
								//MDataIn <= 32'h00000000;
								inPort <= 32'd0;
								clr <= 0;
								//enable[27] <= 0;
								Gra <= 0; 
								Grb <= 0;
								Grc <= 0;
								Rin <= 0;
								Rout <= 0;
								BAout <= 0;
								ReadRAM <= 0;
								WriteRAM <= 0;
								enable[20] <= 1;
								
		end
		Reg_load1a: begin
								//MDataIn <= 32'b0;
								//MD_Read = 0; enable[21] = 0;
								//#10 MD_Read <= 1; enable[21] <= 1;
								////MDataIn <= 32'b0011;
								//#15 MD_Read <= 0; enable[21] <= 0;
								#25 enable[20] <= 1;
								
		end
		Reg_load1b: begin
								//#10 busSelect[21] <= 1; enable[2] <= 1;
								//#15 busSelect[21] <= 0; enable[2] <= 0;
								#25 enable[20] <= 0;
		end
		Reg_load2a: begin
								//MDataIn <= 32'b0110;
								//#10 MD_Read <= 1; enable[21] <= 1;
								//MDataIn <= 32'b0010;
								//#15 MD_Read <= 0; enable[21] <= 0;
								//enable[1] <= 1; ReadRAM <= 1;
		end
		Reg_load2b: begin
								#10 busSelect[21] <= 1; enable[3] <= 1;
								#15 busSelect[21] <= 0; enable[3] <= 0;
		end
		Reg_load3a: begin
								MDataIn <= 32'b0;
								#10 MD_Read <= 1; enable[21] <= 1;
								//MDataIn <= 32'b0;
								#15 MD_Read <= 0; enable[21] <= 0;
		end
		Reg_load3b: begin
								#10 busSelect[21] <= 1; enable[1] <= 1;
								#15 busSelect[21] <= 0; enable[1] <= 0;
		end
		T0: begin
								#10 busSelect[20] <= 1;//PC
								enable[25] <= 1;//MAR
								//enable[27] <= 1;//incPC bit is bit 27
								Control_Signals <= 14;
								enable[18] <= 1;//Zin
								
								#15 busSelect[20] <= 0;
								enable[25] <= 0;//MAR
								//enable[27] <= 0;//incPC bit is bit 27
								Control_Signals <= 0;
								enable[18] <= 0;//Zin
																
		end
		T1: begin
								#10 busSelect[19] <= 1;//zLowOut
								enable[20] <= 1;//pcIn
								enable[21] <= 1;//MDRin
								MD_Read <= 1;//read
								
								//MDataIn <= 32'h0000000010000;//Opcode need to get info into MDR from RAM
								ReadRAM <= 1;
								
								#15 busSelect[19] <= 0;
								busSelect[19] <= 0;
								enable[20] <= 0;
								ReadRAM <= 0;
		end
		T2: begin
							
								#10 enable[21] <= 0; MD_Read <= 0; busSelect[21] <= 1; enable[24] <= 1;
								
								#15 busSelect[21] <= 0; enable[24] <= 0;

		end
		T3: begin
								
								
								
								
								//Gra, Rout and CONIN
								#10 Gra <= 1; busSelect[0] <= 1; enable[27] <= 1;
								#15 Gra <= 0; busSelect[0] <= 0; enable[27] <= 0;
		end
		T4: begin
								
								
								//PC out and Y in
								
								#10 busSelect[20] <=1; enable[19] <= 1;
								#15 busSelect[20] <=0; enable[19] <= 0;
		end
		T5: begin
								
								
								//Cout, ADD, ZIn
								
								#10 busSelect[23] <= 1; enable[18] <= 1;
								#15 busSelect[23] <= 0; enable[18] <= 0;
		end
		T6: begin

								#10 MD_Read <= 1; ReadRAM <= 1; enable[21] <= 1;
								
								#15  ReadRAM <= 0;
		end
		T7: begin

								#10 MD_Read <= 0; enable[21] <= 0; 
								    busSelect[21] <= 1; Gra <= 1; Rin <= 1;
								
								#15 Rin <= 0;
								#15 busSelect[21]<= 0; Gra <= 0;
		end
	endcase
end
endmodule
