module Datapath(
  input wire [31:0] InPort,
  output wire [31:0] OutPort,
  input [31:0] MDatain,
  
);
