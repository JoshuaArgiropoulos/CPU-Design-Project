module ConnectedBus(EncodeIn,
							BusMuxInR0,
							BusMuxInR1,
							BusMuxInR2,
							BusMuxInR3,
							BusMuxInR4,
							BusMuxInR5,
							BusMuxInR6,
							BusMuxInR7,
							BusMuxInR8,
							BusMuxInR9,
							BusMuxInR10,
							BusMuxInR11,
							BusMuxInR12,
							BusMuxInR13,
							BusMuxInR14,
							BusMuxInR15,
							BusMuxInHI,
							BusMuxInLO,
							BusMuxInZHI,
							BusMuxInZLO,
							BusMuxInPc,
							BusMuxInMDR,
							BusMuxInInPort,
							CSignExtended,
							BusMuxOut);
							//EncodeOut
						
						input [31:0] EncodeIn,
							BusMuxInR0,
							BusMuxInR1,
							BusMuxInR2,
							BusMuxInR3,
							BusMuxInR4,
							BusMuxInR5,
							BusMuxInR6,
							BusMuxInR7,
							BusMuxInR8,
							BusMuxInR9,
							BusMuxInR10,
							BusMuxInR11,
							BusMuxInR12,
							BusMuxInR13,
							BusMuxInR14,
							BusMuxInR15,
							BusMuxInHI,
							BusMuxInLO,
							BusMuxInZHI,
							BusMuxInZLO,
							BusMuxInPc,
							BusMuxInMDR,
							BusMuxInInPort,
							CSignExtended;
							//BusMuxOut;

							output [31:0] BusMuxOut;

							wire [4:0] EncodeOut;

Encoder enc_inst(EncodeIn, EncodeOut);
Multiplexer mul_inst(BusMuxInR0,
							BusMuxInR1,
							BusMuxInR2,
							BusMuxInR3,
							BusMuxInR4,
							BusMuxInR5,
							BusMuxInR6,
							BusMuxInR7,
							BusMuxInR8,
							BusMuxInR9,
							BusMuxInR10,
							BusMuxInR11,
							BusMuxInR12,
							BusMuxInR13,
							BusMuxInR14,
							BusMuxInR15,
							BusMuxInHI,
							BusMuxInLO,
							BusMuxInZHI,
							BusMuxInZLO,
							BusMuxInPc,
							BusMuxInMDR,
							BusMuxInInPort,
							CSignExtended,
							BusMuxOut,
							EncodeOut);

endmodule
