module Datapath(
)
